* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 08 Jun 2011 11:13:32 AM EDT


U1  38 37 36 35 34 33 32 31 30 29 1 39 28 27 26 25 24 23 22 21 3 4 5 6 7 8 9 10 11 12 40 2 13 14 15 16 17 18 19 20 PIC18F4620
U2  57 53 55 63 56 50 44 62 52 51 54 45 47 46 43 41 58 44 42 42 44 48 49 61 44 44 60 59 FT232RL
Conn1  42 41 43 44 44 44 CONN USB

.end
